//******************************************************
//COPYRIGHT(c)2016,SouthChina university of technology
//ALL rights reserved.
//IP LIB INDEX :
//IP Name		:
//
//File name		:fbosc2.v
//Module name 	:fbosc2
//Full name		:
//
//Author 		:LeeJT
//Email			:1164880972@qq.com
//Data			:
//Version		:
//
//Abstract		:
//Called by		:Father Module
//
//Modification history
//--------------------------------------------------------
// //
// $LOG$
//
//********************************************************

//********************************************************
//DEFINE MODULE PORT //
//********************************************************
//
module fbosc2 (//INPUT
						clk,
						rst,
					  //OUTPUT
						y1,
						y2
					  );
//********************************************************
//DEFINE PARAMETER //
//********************************************************


//********************************************************
//DEFINE INPUT //
//********************************************************
input clk, rst;
//********************************************************
//DEFINE OUTPUT //
//********************************************************
output y1, y2;
//********************************************************
//OUTPUT ATRIBUTE //
//********************************************************
//REGS
reg y1, y2;

//WIRES



//********************************************************
//MODULE  REGISTERS/WIRES DEFINE //
//********************************************************




//********************************************************
//INSTANCE MODULE //
//********************************************************



//********************************************************
//MAIN CODE //
//********************************************************
always @(posedge clk,posedge rst)
begin 
	if(rst) y2 <=1;
	else y2 <= y1;
end


always @(posedge clk,posedge rst)
begin 
	if(rst) y1 <=0;
	else y1 <= y2;
end

//********************************************************//
endmodule






