library verilog;
use verilog.vl_types.all;
entity fbosc1_vlg_tst is
end fbosc1_vlg_tst;
