library verilog;
use verilog.vl_types.all;
entity fbosc2_vlg_tst is
end fbosc2_vlg_tst;
