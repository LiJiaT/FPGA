//******************************************************
//COPYRIGHT(c)2016,SouthChina university of technology
//ALL rights reserved.
//IP LIB INDEX :
//IP Name		:
//
//File name		:sigdata.v
//Module name 	:sigdata
//Full name		:
//
//Author 		:LeeJT
//Email			:1164880972@qq.com
//Data			:
//Version		:
//
//Abstract		:
//Called by		:Test Module
//
//Modification history
//--------------------------------------------------------
// //
// $LOG$
//
//********************************************************

//********************************************************
//DEFINE MODULE PORT //
//********************************************************
//
`timescale 1ns/1ns
`define halfperiod 50

module sigdata(
					  //INPUT
				ack,
					  //OUTPUT
				rst,
				data,
				sclk
					  );
//********************************************************
//DEFINE PARAMETER //
//********************************************************


//********************************************************
//DEFINE INPUT //
//********************************************************
input ack;
//********************************************************
//DEFINE OUTPUT //
//********************************************************
output rst,sclk;
output [3:0] data;
//********************************************************
//OUTPUT ATRIBUTE //
//********************************************************
//REGS
reg rst,sclk;
reg [3:0] data;

//WIRES



//********************************************************
//MODULE  REGISTERS/WIRES DEFINE //
//********************************************************



//********************************************************
//INSTANCE MODULE //
//********************************************************



//********************************************************
//MAIN CODE //
//********************************************************
initial begin 
	rst =1;
	#10 rst = 0;
	#(`halfperiod*2+3) rst =1;
end

initial begin 
	sclk =0 ;
	data =0;
	#(`halfperiod*1000) $stop;
end


always #(`halfperiod) sclk = ~sclk;

always @(posedge ack)
begin
	#(`halfperiod/2+3) data =data + 1;
end

//********************************************************//
endmodule










