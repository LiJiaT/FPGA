//******************************************************
//COPYRIGHT(c)2016,SouthChina university of technology
//ALL rights reserved.
//IP LIB INDEX :
//IP Name		:
//
//File name		:osc2.v
//Module name 	:osc2
//Full name		:
//
//Author 		:LeeJT
//Email			:1164880972@qq.com
//Data			:
//Version		:
//
//Abstract		:
//Called by		:Father Module
//
//Modification history
//--------------------------------------------------------
// //
// $LOG$
//
//********************************************************

//********************************************************
//DEFINE MODULE PORT //
//********************************************************
//

/*
This is a self-trigger ocilitor generating clock output.
It is a training module for understanding unblock assignment at the begining.
*/


module osc2 (
					  //INPUT
					clk
					  //OUTPUT
						
					  );
//********************************************************
//DEFINE PARAMETER //
//********************************************************


//********************************************************
//DEFINE INPUT //
//********************************************************

//********************************************************
//DEFINE OUTPUT //
//********************************************************
output clk;
//********************************************************
//OUTPUT ATRIBUTE //
//********************************************************
//REGS
reg clk;

//WIRES



//********************************************************
//MODULE  REGISTERS/WIRES DEFINE //
//********************************************************




//********************************************************
//INSTANCE MODULE //
//********************************************************



//********************************************************
//MAIN CODE //
//********************************************************

initial 	
begin
	#10 clk =0;

end

always @(clk) #10 clk <=~clk;

//********************************************************//
endmodule










