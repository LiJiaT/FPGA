module CPU (data,rst,clk,opcode,ir_addr,opcode,ir_addr,rd,wr,halt,dataout,addr);
input [7:0] data;
input rst,clk;
input [2:0] opcode, ir_addr;

output [2:0] opcode, ir_addr

endmodule