library verilog;
use verilog.vl_types.all;
entity EEPROM_I2CWR is
    generic(
        IDLE            : vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        Ready           : vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        Write_start     : vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        Ctrl_write      : vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        Addr_write      : vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        Data_write      : vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        Read_start      : vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        Ctrl_read       : vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        Data_read       : vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        Stop            : vl_logic_vector(0 to 10) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        Ackn            : vl_logic_vector(0 to 10) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        sh8out_bit7     : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        sh8out_bit6     : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        sh8out_bit5     : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        sh8out_bit4     : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        sh8out_bit3     : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        sh8out_bit2     : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        sh8out_bit1     : vl_logic_vector(0 to 8) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        sh8out_bit0     : vl_logic_vector(0 to 8) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        sh8out_end      : vl_logic_vector(0 to 8) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        sh8in_begin     : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        sh8in_bit7      : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        sh8in_bit6      : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        sh8in_bit5      : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        sh8in_bit4      : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        sh8in_bit3      : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        sh8in_bit2      : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        sh8in_bit1      : vl_logic_vector(0 to 9) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        sh8in_bit0      : vl_logic_vector(0 to 9) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        sh8in_end       : vl_logic_vector(0 to 9) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        head_begin      : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        head_bit        : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        head_end        : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        stop_begin      : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        stop_bit        : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        stop_end        : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        YES             : vl_logic := Hi1;
        NO              : vl_logic := Hi0
    );
    port(
        rst             : in     vl_logic;
        CLK             : in     vl_logic;
        WR              : in     vl_logic;
        RD              : in     vl_logic;
        ADDR            : in     vl_logic_vector(10 downto 0);
        SDA             : inout  vl_logic;
        DATA            : inout  vl_logic_vector(7 downto 0);
        SCL             : out    vl_logic;
        ACK             : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of IDLE : constant is 1;
    attribute mti_svvh_generic_type of Ready : constant is 1;
    attribute mti_svvh_generic_type of Write_start : constant is 1;
    attribute mti_svvh_generic_type of Ctrl_write : constant is 1;
    attribute mti_svvh_generic_type of Addr_write : constant is 1;
    attribute mti_svvh_generic_type of Data_write : constant is 1;
    attribute mti_svvh_generic_type of Read_start : constant is 1;
    attribute mti_svvh_generic_type of Ctrl_read : constant is 1;
    attribute mti_svvh_generic_type of Data_read : constant is 1;
    attribute mti_svvh_generic_type of Stop : constant is 1;
    attribute mti_svvh_generic_type of Ackn : constant is 1;
    attribute mti_svvh_generic_type of sh8out_bit7 : constant is 1;
    attribute mti_svvh_generic_type of sh8out_bit6 : constant is 1;
    attribute mti_svvh_generic_type of sh8out_bit5 : constant is 1;
    attribute mti_svvh_generic_type of sh8out_bit4 : constant is 1;
    attribute mti_svvh_generic_type of sh8out_bit3 : constant is 1;
    attribute mti_svvh_generic_type of sh8out_bit2 : constant is 1;
    attribute mti_svvh_generic_type of sh8out_bit1 : constant is 1;
    attribute mti_svvh_generic_type of sh8out_bit0 : constant is 1;
    attribute mti_svvh_generic_type of sh8out_end : constant is 1;
    attribute mti_svvh_generic_type of sh8in_begin : constant is 1;
    attribute mti_svvh_generic_type of sh8in_bit7 : constant is 1;
    attribute mti_svvh_generic_type of sh8in_bit6 : constant is 1;
    attribute mti_svvh_generic_type of sh8in_bit5 : constant is 1;
    attribute mti_svvh_generic_type of sh8in_bit4 : constant is 1;
    attribute mti_svvh_generic_type of sh8in_bit3 : constant is 1;
    attribute mti_svvh_generic_type of sh8in_bit2 : constant is 1;
    attribute mti_svvh_generic_type of sh8in_bit1 : constant is 1;
    attribute mti_svvh_generic_type of sh8in_bit0 : constant is 1;
    attribute mti_svvh_generic_type of sh8in_end : constant is 1;
    attribute mti_svvh_generic_type of head_begin : constant is 1;
    attribute mti_svvh_generic_type of head_bit : constant is 1;
    attribute mti_svvh_generic_type of head_end : constant is 1;
    attribute mti_svvh_generic_type of stop_begin : constant is 1;
    attribute mti_svvh_generic_type of stop_bit : constant is 1;
    attribute mti_svvh_generic_type of stop_end : constant is 1;
    attribute mti_svvh_generic_type of YES : constant is 1;
    attribute mti_svvh_generic_type of NO : constant is 1;
end EEPROM_I2CWR;
