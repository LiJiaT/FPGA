library verilog;
use verilog.vl_types.all;
entity EEPROM_I2CWR_vlg_tst is
end EEPROM_I2CWR_vlg_tst;
